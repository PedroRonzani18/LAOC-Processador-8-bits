library verilog;
use verilog.vl_types.all;
entity BancoDeRegistradores_simulacao is
end BancoDeRegistradores_simulacao;
