library verilog;
use verilog.vl_types.all;
entity ULA_simulacao is
end ULA_simulacao;
