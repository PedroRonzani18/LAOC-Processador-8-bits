library verilog;
use verilog.vl_types.all;
entity MenoriaInstrucao_simulacao is
end MenoriaInstrucao_simulacao;
