library verilog;
use verilog.vl_types.all;
entity \AND\ is
    port(
        Entrada1        : in     vl_logic;
        Entrada2        : in     vl_logic;
        Resultado       : out    vl_logic
    );
end \AND\;
