library verilog;
use verilog.vl_types.all;
entity MUX3_3_simulacao is
end MUX3_3_simulacao;
