library verilog;
use verilog.vl_types.all;
entity PC_simulacao is
end PC_simulacao;
