library verilog;
use verilog.vl_types.all;
entity armazenaEstados is
end armazenaEstados;
