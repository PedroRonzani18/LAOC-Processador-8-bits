library verilog;
use verilog.vl_types.all;
entity ExtensorDeSinal_simulacao is
end ExtensorDeSinal_simulacao;
