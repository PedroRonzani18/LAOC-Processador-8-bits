library verilog;
use verilog.vl_types.all;
entity MenoriaDados_simulacao is
end MenoriaDados_simulacao;
