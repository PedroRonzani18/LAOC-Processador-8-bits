library verilog;
use verilog.vl_types.all;
entity MUX3_8_simulacao is
end MUX3_8_simulacao;
