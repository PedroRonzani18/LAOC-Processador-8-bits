library verilog;
use verilog.vl_types.all;
entity Somador_simulacao is
end Somador_simulacao;
