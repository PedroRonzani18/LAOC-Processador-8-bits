library verilog;
use verilog.vl_types.all;
entity MUX2_8_simulacao is
end MUX2_8_simulacao;
