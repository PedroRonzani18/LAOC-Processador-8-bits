library verilog;
use verilog.vl_types.all;
entity UnidadeControle_simulacao is
end UnidadeControle_simulacao;
