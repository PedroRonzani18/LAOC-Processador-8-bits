library verilog;
use verilog.vl_types.all;
entity AND_simulacao is
end AND_simulacao;
