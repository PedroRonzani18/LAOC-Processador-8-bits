library verilog;
use verilog.vl_types.all;
entity MUX2_3_simulacao is
end MUX2_3_simulacao;
